//-----------------------$finish()----------------------------//
task finish();
#(run_time)
$display("!!!!!!!!!!!!!!!!!!!!!!!END OF TB!!!!!!!!!!!!!!!!!!!!!!!!!!!!");
$finish(1);
endtask
//-------------------------------------------------------------//